module company

import freeflowuniverse.baobab.modelbase
// import freeflowuniverse.baobab.modelactors.finance
// import freeflowuniverse.baobab.modelglobal.country
import freeflowuniverse.crystallib.timetools { time_from_string }
import freeflowuniverse.crystallib.params { Tags ParamsFilter}
import time

// budget_item
// This file deals with the budget item base and...


