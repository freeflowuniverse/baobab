module modelglobal

import time

[heap]
struct DBGLBase {
pub mut:
	dbgl &DBGLData
}
