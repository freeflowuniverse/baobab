module processor

